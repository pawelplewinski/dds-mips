library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity mips32sys is 
    generic (
        PGM_FILE 	: string   := "no.file";
        IA_LEN      : natural  :=  9;
		DA_LEN      : natural  :=  6;
        GPIO_LEN    : natural  :=  8
    );
    port(
        clk         : in  std_logic;
        resetn      : in  std_logic
    );
end entity mips32sys;
    
architecture gut_struct of mips32sys is

    ---------------
    -- MIPS core --
    ---------------
    component mips32core is
    generic(
        IA_LEN    : natural  :=  9
    );
    port(
        ibus_data_inp   : in  std_logic_vector(31 downto 0);
        ibus_addr_out   : out std_logic_vector(31 downto 0);
        
        dbus_addr_out   : out std_logic_vector(31 downto 0);
        dbus_data_inp   : in  std_logic_vector(31 downto 0);
        dbus_data_out   : out std_logic_vector(31 downto 0);
        dbus_wren_out   : out std_logic;
        
        clk             : in std_logic;
        resetn          : in std_logic
    );
    end component mips32core;

    ------------
    -- memory --
    ------------
    component mem32 is
    generic(
        PGM_FILE 	: string  := "no.file";
        ADDR_LENGTH : natural :=  9
    );
    port(
        -- COM bus interface
        bus_addr_inp    : in  std_logic_vector(31 downto 0);
        bus_data_inp    : in  std_logic_vector(31 downto 0);
        bus_data_out    : out std_logic_vector(31 downto 0);
        bus_wren_inp    : in  std_logic;                                        -- '1' -> enable write ; '0' -> disable write
          
        clk             : in std_logic;
        resetn          : in std_logic
    );
    end component mem32;
    
    -- Use the different flavours of the memory component
    for imem : mem32 use entity work.mem32(ibehav);
    for dmem : mem32 use entity work.mem32(dbehav);
  
    ---------------------------------------
    --------------- Signals ---------------
    ---------------------------------------
    
    -- bus signals for COM with RAM components from the master PoV (core -> I/O) 
    -- imem(iram):
    --signal iram_d_i   : std_logic_vector(SYS_32-1 downto 0);        -- [obsolete] holds new instr data for imem
    signal iram_data_inp    : std_logic_vector(31 downto 0);        -- holds new instr from imem
    signal iram_addr_out    : std_logic_vector(31 downto 0);        -- holds new instr addr for imem
    --signal iram_we_o  : std_logic;                                  -- [obsolete] holds the write enable signal from core->imem
    -- dmem(dram):
    signal dram_data_inp    : std_logic_vector(31 downto 0);
    signal dram_addr_out    : std_logic_vector(31 downto 0);
    signal dram_data_out    : std_logic_vector(31 downto 0);
    signal dram_wren_out    : std_logic;
    
begin

    -- Connect MIPS core
    cpu : entity work.mips32core(behavior)
        generic map(
            IA_LEN          => IA_LEN
        )
        port map(
            ibus_data_inp   => iram_data_inp,
            ibus_addr_out   => iram_addr_out,

            dbus_data_inp   => dram_data_inp,
            dbus_addr_out   => dram_addr_out,
            dbus_data_out   => dram_data_out,
            dbus_wren_out   => dram_wren_out,

            clk             => clk,
            resetn          => resetn
        );

    -- Connect instruction memory
    imem : mem32
        generic map(
            PGM_FILE 	    => PGM_FILE,
            ADDR_LENGTH     => IA_LEN
        )
        port map(
            bus_wren_inp    => '0',             -- only read imem memory
            bus_addr_inp    => iram_addr_out,
            bus_data_inp    => (others => 'Z'), -- no write data 
            bus_data_out    => iram_data_inp,
           
            clk             => clk,
            resetn          => resetn
        );

    -- Connect data memory            
    dmem : mem32
        generic map(
            ADDR_LENGTH     => DA_LEN
        )
        port map(
            bus_wren_inp    => dram_wren_out,
            bus_addr_inp    => dram_addr_out,
            bus_data_inp    => dram_data_out,
            bus_data_out    => dram_data_inp,

            clk             => clk,
            resetn          => resetn
        );

end architecture gut_struct;

    
architecture dut_struct of mips32sys is

    ---------------
    -- MIPS core --
    ---------------
    component mips32core is
    generic(
        IA_LEN    : natural  :=  9
    );
    port(
        ibus_data_inp   : in  std_logic_vector(31 downto 0);
        ibus_addr_out   : out std_logic_vector(31 downto 0);
        
        dbus_addr_out   : out std_logic_vector(31 downto 0);
        dbus_data_inp   : in  std_logic_vector(31 downto 0);
        dbus_data_out   : out std_logic_vector(31 downto 0);
        dbus_wren_out   : out std_logic;
        
        clk             : in std_logic;
        resetn          : in std_logic
    );
    end component mips32core;

    ------------
    -- memory --
    ------------
    component mem32 is
    generic(
        PGM_FILE 	: string := "no.file";
        ADDR_LENGTH : natural  :=  9
    );
    port(
        -- COM bus interface
        bus_addr_inp    : in  std_logic_vector(31 downto 0);
        bus_data_inp    : in  std_logic_vector(31 downto 0);
        bus_data_out    : out std_logic_vector(31 downto 0);
        bus_wren_inp    : in  std_logic;                                        -- '1' -> enable write ; '0' -> disable write
          
        clk             : in std_logic;
        resetn          : in std_logic
    );
    end component mem32;
    
    -- Use the different flavours of the memory component
    for imem : mem32 use entity work.mem32(ibehav);
    for dmem : mem32 use entity work.mem32(dbehav);
  
    ---------------------------------------
    --------------- Signals ---------------
    ---------------------------------------
    
    -- bus signals for COM with RAM components from the master PoV (core -> I/O) 
    -- imem(iram):
    --signal iram_d_i   : std_logic_vector(SYS_32-1 downto 0);        -- [obsolete] holds new instr data for imem
    signal iram_data_inp    : std_logic_vector(31 downto 0);        -- holds new instr from imem
    signal iram_addr_out    : std_logic_vector(31 downto 0);        -- holds new instr addr for imem
    --signal iram_we_o  : std_logic;                                  -- [obsolete] holds the write enable signal from core->imem
    -- dmem(dram):
    signal dram_data_inp    : std_logic_vector(31 downto 0);
    signal dram_addr_out    : std_logic_vector(31 downto 0);
    signal dram_data_out    : std_logic_vector(31 downto 0);
    signal dram_wren_out    : std_logic;
    
begin

    -- Connect MIPS core
    cpu : entity work.mips32core(structural)
        generic map(
            IA_LEN          => IA_LEN
        )
        port map(
            ibus_data_inp   => iram_data_inp,
            ibus_addr_out   => iram_addr_out,

            dbus_data_inp   => dram_data_inp,
            dbus_addr_out   => dram_addr_out,
            dbus_data_out   => dram_data_out,
            dbus_wren_out   => dram_wren_out,

            clk             => clk,
            resetn          => resetn
        );

    -- Connect instruction memory
    imem : mem32
        generic map(
            PGM_FILE 	    => PGM_FILE,
            ADDR_LENGTH     => IA_LEN
        )
        port map(
            bus_wren_inp    => '0',             -- only read imem memory
            bus_addr_inp    => iram_addr_out,
            bus_data_inp    => (others => 'Z'), -- no write data 
            bus_data_out    => iram_data_inp,
           
            clk             => clk,
            resetn          => resetn
        );

    -- Connect data memory            
    dmem : mem32
        generic map(
            ADDR_LENGTH     => DA_LEN
        )
        port map(
            bus_wren_inp    => dram_wren_out,
            bus_addr_inp    => dram_addr_out,
            bus_data_inp    => dram_data_out,
            bus_data_out    => dram_data_inp,

            clk             => clk,
            resetn          => resetn
        );

end architecture dut_struct;